#!/usr/bin/python3
import sys
import os
import colorama
from colorama import Fore, Style

if sys.argv[0] != "./ckt":
    print("Comando no valido.")
    exit(0)

def printHelp():
    print("Chikatana Command Line:")

if len(sys.argv) == 1:
    printHelp()
    exit(0)

if sys.argv[1] == "init":
    os.system("docker-compose up -d")
    exit(0)

if sys.argv[1] == "up":
    os.system("docker-compose up -d")
    exit(0)

if sys.argv[1] == "down":
    os.system("docker-compose down")
    exit(0)

if sys.argv[1] == "ps":
    print(Fore.CYAN + "Monstando contenedores ..." + Style.RESET_ALL)
    os.system("docker-compose ps")
    exit(0)

if sys.argv[1] == "restart":
    os.system("docker-compose down && docker-compose up -d")
    exit(0)




###################################################################################
#                                                                                 #
#                                 DB COMMANDS                                #
#                                                                                 #
###################################################################################

if sys.argv[1] == "db":
    if len(sys.argv) == 2:
        os.system("docker-compose exec -u www-data db mysql -u magento -p magento")
        exit(0)
    elif len(sys.argv) >= 3:
        if sys.argv[2] == "clean":
            print("Eliminando y creando base de datos")
            query = """
                DROP DATABASE magento;
                CREATE DATABASE magento;
                """
            os.system("docker-compose exec -u www-data db mysql -u magento -p -e \"" + query + "\"")
            print("Listo.")
            exit(0)
        elif sys.argv[2] == "fix":
            hostname = 'https://magento.ckt/'
            print("Comenzara el fix")
            query = """
                UPDATE core_config_data SET value='%s' WHERE path='web/unsecure/base_url';
                UPDATE core_config_data SET value='%s' WHERE path='web/secure/base_url';
                UPDATE core_config_data SET value='%s' WHERE path='web/unsecure/base_link_url';
                UPDATE core_config_data SET value='%s' WHERE path='web/secure/base_link_url';
                """ % (hostname, hostname, hostname, hostname)
            os.system("docker-compose exec -u root db mysql -u magento -p magento -e \"" + query + "\"")
            print("Listo.")
            exit(0)

        # Mensaje para indicar que el comando no fue encontrado
        print("El comando esta incorrecto")
    else:
        # Mensaje para indicar que el comando no se puede ejecutar
        print("El comando esta incompleto")
    exit(0)




###################################################################################
#                                                                                 #
#                                 MAGENTO COMMANDS                                #
#                                                                                 #
###################################################################################

if sys.argv[1] == "adobe":
    if len(sys.argv) == 2:
        os.system("docker-compose exec -u magento2 web bash")
        exit(0)
    elif len(sys.argv) >= 3:
        if sys.argv[2] == "composer":
            os.system("docker-compose exec -u magento2 web composer install")
            exit(0)
        elif sys.argv[2] == "upgrade":
            os.system("docker-compose exec -u magento2 web php bin/magento setup:upgrade")
            exit(0)
        elif sys.argv[2] == "reindex":
            os.system("docker-compose exec -u magento2 web php bin/magento indexer:reindex")
            exit(0)



        ###########################################################################
        #                             CACHE COMMANDS                              #
        ###########################################################################

        elif sys.argv[2] == "cache":
            if len(sys.argv) == 3:
                print(Fore.CYAN + "Limpiando Cache ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento cache:clean")
                print(Fore.CYAN + "Hecho." + Style.RESET_ALL)
                exit(0)
            elif sys.argv[3] == "status":
                os.system("docker-compose exec -u magento2 web php bin/magento cache:status")
                exit(0)
            elif sys.argv[3] == "enable":
                print(Fore.BLUE + "Enable Cahe ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento cache:enable")
                print(Fore.BLUE + "Disable Cahe Modules ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento cache:disable collections eav full_page layout")
                print(Fore.GREEN + "Hecho." + Style.RESET_ALL)
                exit(0)
            elif sys.argv[3] == "disable":
                print(Fore.BLUE + "Disable Cahe ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento cache:disable")
                print(Fore.GREEN + "Hecho." + Style.RESET_ALL)
                exit(0)
            elif sys.argv[3] == "clear":
                print(Fore.BLUE + "Clear Cahe ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento cache:clean")
                # print(Fore.BLUE + "Cambiando permisos ..." + Style.RESET_ALL)
                # os.system("docker-compose exec -u magento2 web chown -R magento2:magento2 generated pub var")
                print(Fore.GREEN + "Hecho." + Style.RESET_ALL)
                exit(0)
            else:
                print("El comando de magento esta incompleto")



        ###########################################################################
        #                             RESET COMMANDS                              #
        ###########################################################################

        elif sys.argv[2] == "reset":
            print(Fore.CYAN + "Bajando contenedores..." + Style.RESET_ALL)
            os.system("docker-compose down")
            print(Fore.CYAN + "Eliminando archivos cache y estaticos..." + Style.RESET_ALL)
            os.system("rm -rf generated/* pub/static/*")
            print(Fore.CYAN + "Levantando contenedores..." + Style.RESET_ALL)
            os.system("docker-compose up -d")
            print(Fore.CYAN + "Actualizando Magento..." + Style.RESET_ALL)
            os.system("docker-compose exec -u magento2 web php bin/magento setup:upgrade")
            print(Fore.CYAN + "Actilizando cache de Magento..." + Style.RESET_ALL)
            os.system("docker-compose exec -u magento2 web php bin/magento cache:clean")
            print(Fore.CYAN + "Comando finalizado." + Style.RESET_ALL)
            exit(0)



        ###########################################################################
        #                         TEMPLATE HINTS COMMANDS                         #
        ###########################################################################

        elif sys.argv[2] == "template-hints":
            if len(sys.argv) == 4 and sys.argv[3] == "enable":
                print(Fore.BLUE + "Enable template hints ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento dev:template-hints:enable")
            else:
                print(Fore.BLUE + "Disable template hints ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento dev:template-hints:disable")

            print(Fore.BLUE + "Clear Cahe ..." + Style.RESET_ALL)
            os.system("docker-compose exec -u magento2 web php bin/magento cache:clean")
            print(Fore.GREEN + "Hecho." + Style.RESET_ALL)
            exit(0)



        ###########################################################################
        #                             STYLES COMMANDS                             #
        ###########################################################################

        elif sys.argv[2] == "styles":
            print(Fore.BLUE + "Compilando Estilos ..." + Style.RESET_ALL)
            os.system("docker-compose exec -u magento2 web grunt clean exec:biz less:biz;")
            print(Fore.BLUE + "Borrando Cahe ..." + Style.RESET_ALL)
            os.system("docker-compose exec -u magento2 web php bin/magento cache:clean")
            print(Fore.GREEN + "Hecho." + Style.RESET_ALL)
            exit(0)



        ###########################################################################
        #                             STYLES COMMANDS                             #
        ###########################################################################

        elif sys.argv[2] == "static-content":
            print(Fore.CYAN + "Deploy static content ..." + Style.RESET_ALL)
            os.system("docker-compose exec -u magento2 web php bin/magento setup:static-content:deploy es_MX -f")
            print(Fore.CYAN + "Hecho." + Style.RESET_ALL)
            exit(0)


        ###########################################################################
        #                             OTHERS COMMANDS                             #
        ###########################################################################

        elif sys.argv[2] == "create":
            if  sys.argv[3] == "admin-user":
                print(Fore.BLUE + "Creando Palomino admin ..." + Style.RESET_ALL)
                os.system("docker-compose exec -u magento2 web php bin/magento admin:user:create --admin-user='palomino' --admin-password='Law200110513' --admin-email='palomino@wolfsellers.com' --admin-firstname='palomino' --admin-lastname='palomino'")
            else:
                print("No se encontro el commando a ejecutar.")
            exit(0)


        # Mensaje para indicar que el comando no fue encontrado
        print("El comando docker no encontrado")
    else:
        # Mensaje para indicar que el comando no se puede ejecutar
        print("El comando de magento esta incompleto")
    exit(0)
